`include "uvm_macros.svh"

package apb_pkg;

    import uvm_pkg::*;
    
    `include "apb_data_item.sv"
    `include "apb_seqlib.sv"
    // `include "apb_master_driver.sv"

endpackage